CLK28MPLL_DE2_115_inst : CLK28MPLL_DE2_115 PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig,
		c1	 => c1_sig
	);
